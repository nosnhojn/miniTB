module dut();
endmodule
