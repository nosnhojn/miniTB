module dut;
reg a;
endmodule
